
  localparam CLK_FREQ   = 50000000;

  localparam LED_FREQ_STEPS = 10;
  localparam LED_MAX_FREQ   = 110;
  localparam LED_MIN_FREQ   = 10;
  localparam LED_SCALE_DIV  = 1;
  localparam LED_INIT_STEP  = 4;

  localparam TICK_FREQ_STEPS = 4;
  localparam TICK_MAX_FREQ   = 50;
  localparam TICK_MIN_FREQ   = 1;
  localparam TICK_SCALE_DIV  = 10;
  localparam TICK_INIT_STEP  = 2;

  localparam NUM_SYNC   = 3;
  localparam DEBOUNCE   = 16;
  localparam BTN_ACTIVE = 0;
  localparam LED_WIDTH  = 8;
